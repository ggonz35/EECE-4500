library ieee;
library vga;
library ads;
library algor;



