library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use std.textio.all;

use work.ads.all;
use work.vga.all;

entity mandelbrot is
	port(
		clk_50 			: in std_logic;
		vga_vs 			: out std_logic;			
		vga_hs 			: out std_logic;
		vga_r 			: out std_logic(0 to 3);
		vga_g 			: out std_logic(0 to 3);
		vga_b 			: out std_logic(0 to 3)
		
	);
end mandelbrot;

architecture steve of mandelbrot is
	
	signal vga_clk		: std_logic_vector (4 downto 0);
	signal rst			: std_logic;
	signal point_out	: coordinate;
	signal p_val_out	: boolean;
	signal vs_out 		: std_logic;
	signal hs_out 		: std_logic;
	signal r_out		: std_logic_vector(0 to 3);
	signal g_out		: std_logic_vector(0 to 3);
	signal b_out		: std_logic_vector(0 to 3);
	signal a_set		: std_logic := '0';
	signal l_set		: std_logic;

begin
    -- Add your VGA configuration and color map setup here
	 
	pll :entity vga_pll 
	
		port map (
		
		arset				<= a_set,
		in_clk			<= clk_50,
		
		vga_clk 			<= c0,
		l_set 			<= locked
		
	);
	
	
	vga:entity vga_fsm
	
		  port map(
		  
		  vga_clock		<= vga_clk,
        reset			<= rst,

		  point_out		<=	point,
		  p_val_out		<= point_valid,

		  vs_out			<= h_sync,
		  hs_out			<= v_sync
		
	);
	
	
	 

end architecture steve;
