* Main Circuit - Includes subcircuit definitions and the ring oscillator with NAND gate

* Define parameters for process variations
.param tplv = 1.0
.param tpwv = 1.0
.param tnln = 1.0
.param tnwn = 1.0
.param tpotv = 1.0
.param tnotv = 1.0

* Include the subcircuit for the inverter
.include inverter.cir

* Include the subcircuit for the NAND gate
.include nand.cir

* Define the ring oscillator with 12 inverters
X1 in1 out1 inverter L=tplv*130n W=tpwv*130n
X2 out1 in2 inverter L=tplv*130n W=tpwv*130n
X3 in2 out2 inverter L=tplv*130n W=tpwv*130n
X4 out2 in3 inverter L=tplv*130n W=tpwv*130n
X5 in3 out3 inverter L=tplv*130n W=tpwv*130n
X6 out3 in4 inverter L=tplv*130n W=tpwv*130n
X7 in4 out4 inverter L=tplv*130n W=tpwv*130n
X8 out4 in5 inverter L=tplv*130n W=tpwv*130n
X9 in5 out5 inverter L=tplv*130n W=tpwv*130n
X10 out5 in6 inverter L=tplv*130n W=tpwv*130n
X11 in6 out6 inverter L=tplv*130n W=tpwv*130n
X12 out6 in1 inverter L=tplv*130n W=tpwv*130n

* Define the enable signal
Venable enable 0 PULSE(0 1 0 1n 1n 0.01n 0.02n 100n) DC 0

* Connect the NAND gate to the ring oscillator with an enable signal
X13 in1 enable out1_nand nand
X14 out1_nand in2 out1_nand nand
